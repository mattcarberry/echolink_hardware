-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Saturday, July 16, 2016 15:06:18 Pacific Daylight Time

